`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/04/2015 12:44:37 AM
// Design Name: 
// Module Name: bitcrusher
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bitcrusher(
    input clock,
    input reset,
    input start,
    input [11:0] incoming_sample,
    output [11:0] modified_sample,
    output done
    );
    
    
    
    
    
endmodule
