module soundproc(input micsound, output success);



endmodule
