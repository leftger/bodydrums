`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/25/2015 01:11:03 AM
// Design Name: 
// Module Name: triangle
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module triangle(
    input [10:0] p_one_x, p_two_x, p_three_x,
    input [10:0] hcount,
    input [9:0] p_one_y, p_two_y, p_three_y,
    input [9:0] vcount,
    output [23:0] pixel
    );
endmodule
