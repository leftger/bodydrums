module soundproc(input micsound, output success);

assign success = 1;

endmodule
